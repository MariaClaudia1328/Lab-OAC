//------------------------------------
// Colocar todos os módulos do processador aqui
//------------------------------------

module processador-uniciclo;



endmodule 